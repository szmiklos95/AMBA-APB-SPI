`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:30:18 05/22/2018 
// Design Name: 
// Module Name:    APB_interface 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module APB_interface(
		input PCLK,
		input PRESETn,
		input [15:0] data_in,
		output [15:0] data_out,
		input [15:0] PWDATA,
		output [15:0] PRDATA
    );


endmodule
